LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

ENTITY DECODIFICADOR_MSG2 IS
	PORT(HABILITACION: IN STD_LOGIC;
	ANODO: OUT STD_LOGIC_VECTOR(6 DOWNTO 0));
END DECODIFICADOR_MSG2;

ARCHITECTURE SOL OF DECODIFICADOR_MSG2 IS
BEGIN
	PROCESS(HABILITACION)
	BEGIN
		CASE HABILITACION IS
			WHEN '1' => ANODO<="1110110";
			WHEN others => ANODO<="0000000";
		END CASE;
	END PROCESS;
END SOL;