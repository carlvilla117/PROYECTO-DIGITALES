LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

ENTITY COMPARADOR IS
	PORT ( A,B: IN STD_LOGIC_VECTOR(3 DOWNTO 0);
		 MY,IG,MN: OUT STD_LOGIC);
END COMPARADOR;

ARCHITECTURE SOL OF COMPARADOR IS
BEGIN
	MY <= '1' WHEN (A>B) ELSE '0';
	IG <= '1' WHEN (A=B) ELSE '0';
	MN <= '1' WHEN (A<B) ELSE '0';
END SOL;