LIBRARY IEEE;
USE ieee.std_logic_1164.all;

ENTITY OR_10 IS
PORT (x : IN STD_LOGIC_VECTOR(9 TO 0);
		f : OUT STD_LOGIC);
END OR_10;

ARCHITECTURE SOL OF OR_10 IS
SIGNAL tmp : STD_LOGIC_VECTOR(9 TO 0);
BEGIN
tmp <= (OTHERS => '0');
f <= '0' WHEN x = tmp ELSE '1';
END SOL;